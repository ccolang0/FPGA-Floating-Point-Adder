`timescale 1ns / 1ps

module FPA_Top(

    );
endmodule
