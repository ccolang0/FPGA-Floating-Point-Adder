`timescale 1ns / 1ps

module FPA_Controller(

    );
endmodule
